module colorconvert(//input data,
							output logic[7:0]red,
							output logic[7:0]green,
							output logic[7:0]blue);
always_comb
begin :RGB_Display
				/*if(data==1)
				begin	
					red=2'h3f;
					green=2'h00;
					blue=2'h3f;
				end
				else
				begin	
					red=2'h3f;
					green=2'h00;
					blue=2'h3f;
				end*/
				
end
endmodule
				